module hello;
  initial begin
    $display("Hello, Verilog! im test the verilog languages so what this can do ");
    $finish;
  end
endmodule
// test 
// test 